// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Sat Mar 25 22:07:02 2017"

module InstructionFetch(
	CW
);


output wire	[55:0] CW;

wire	[55:0] CW_ALTERA_SYNTHESIZED;






assign	CW = CW_ALTERA_SYNTHESIZED;
assign	CW_ALTERA_SYNTHESIZED[53] = 0;
assign	CW_ALTERA_SYNTHESIZED[52] = 0;
assign	CW_ALTERA_SYNTHESIZED[51] = 0;
assign	CW_ALTERA_SYNTHESIZED[50] = 0;
assign	CW_ALTERA_SYNTHESIZED[49] = 0;
assign	CW_ALTERA_SYNTHESIZED[48] = 0;
assign	CW_ALTERA_SYNTHESIZED[47] = 0;
assign	CW_ALTERA_SYNTHESIZED[46] = 0;
assign	CW_ALTERA_SYNTHESIZED[45] = 0;
assign	CW_ALTERA_SYNTHESIZED[44] = 0;
assign	CW_ALTERA_SYNTHESIZED[43] = 0;
assign	CW_ALTERA_SYNTHESIZED[42] = 0;
assign	CW_ALTERA_SYNTHESIZED[41] = 0;
assign	CW_ALTERA_SYNTHESIZED[40] = 0;
assign	CW_ALTERA_SYNTHESIZED[39] = 0;
assign	CW_ALTERA_SYNTHESIZED[38] = 0;
assign	CW_ALTERA_SYNTHESIZED[37] = 0;
assign	CW_ALTERA_SYNTHESIZED[36] = 0;
assign	CW_ALTERA_SYNTHESIZED[35] = 0;
assign	CW_ALTERA_SYNTHESIZED[34] = 0;
assign	CW_ALTERA_SYNTHESIZED[33] = 0;
assign	CW_ALTERA_SYNTHESIZED[32] = 0;
assign	CW_ALTERA_SYNTHESIZED[31] = 0;
assign	CW_ALTERA_SYNTHESIZED[30] = 0;
assign	CW_ALTERA_SYNTHESIZED[29] = 0;
assign	CW_ALTERA_SYNTHESIZED[28] = 0;
assign	CW_ALTERA_SYNTHESIZED[27] = 0;
assign	CW_ALTERA_SYNTHESIZED[26] = 0;
assign	CW_ALTERA_SYNTHESIZED[25] = 0;
assign	CW_ALTERA_SYNTHESIZED[24] = 0;
assign	CW_ALTERA_SYNTHESIZED[23] = 0;
assign	CW_ALTERA_SYNTHESIZED[22] = 0;
assign	CW_ALTERA_SYNTHESIZED[21] = 0;
assign	CW_ALTERA_SYNTHESIZED[20] = 0;
assign	CW_ALTERA_SYNTHESIZED[19] = 0;
assign	CW_ALTERA_SYNTHESIZED[18] = 0;
assign	CW_ALTERA_SYNTHESIZED[17] = 0;
assign	CW_ALTERA_SYNTHESIZED[16] = 0;
assign	CW_ALTERA_SYNTHESIZED[15] = 0;
assign	CW_ALTERA_SYNTHESIZED[14] = 0;
assign	CW_ALTERA_SYNTHESIZED[13] = 0;
assign	CW_ALTERA_SYNTHESIZED[12] = 0;
assign	CW_ALTERA_SYNTHESIZED[11] = 0;
assign	CW_ALTERA_SYNTHESIZED[10] = 0;
assign	CW_ALTERA_SYNTHESIZED[9] = 0;
assign	CW_ALTERA_SYNTHESIZED[7] = 0;
assign	CW_ALTERA_SYNTHESIZED[6] = 0;
assign	CW_ALTERA_SYNTHESIZED[5] = 0;
assign	CW_ALTERA_SYNTHESIZED[4] = 0;
assign	CW_ALTERA_SYNTHESIZED[2] = 0;
assign	CW_ALTERA_SYNTHESIZED[0] = 0;
assign	CW_ALTERA_SYNTHESIZED[55] = 0;
assign	CW_ALTERA_SYNTHESIZED[3] = 1;
assign	CW_ALTERA_SYNTHESIZED[54] = 1;
assign	CW_ALTERA_SYNTHESIZED[1] = 1;
assign	CW_ALTERA_SYNTHESIZED[8] = 1;

endmodule
