// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Tue Mar 28 23:10:02 2017"

module Ex0_Select(
	IR_in,
	S1,
	S0
);


input wire	[15:0] IR_in;
output wire	S1;
output wire	S0;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;




assign	SYNTHESIZED_WIRE_4 = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_6 | IR_in[10];

assign	S0 = SYNTHESIZED_WIRE_2 | IR_in[13];

assign	SYNTHESIZED_WIRE_0 =  ~IR_in[9];

assign	SYNTHESIZED_WIRE_2 = IR_in[12] & SYNTHESIZED_WIRE_6;

assign	S1 = SYNTHESIZED_WIRE_4 & IR_in[12] & SYNTHESIZED_WIRE_5;

assign	SYNTHESIZED_WIRE_5 =  ~IR_in[13];

assign	SYNTHESIZED_WIRE_6 =  ~IR_in[11];


endmodule
