// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Tue Mar 07 00:51:41 2017"

module \2to4Decoder_2Inputs (
	A,
	B,
	m0,
	m1,
	m2,
	m3
);


input wire	A;
input wire	B;
output wire	m0;
output wire	m1;
output wire	m2;
output wire	m3;

wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;




assign	m0 = SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_5;

assign	m1 = B & SYNTHESIZED_WIRE_5;

assign	m2 = SYNTHESIZED_WIRE_4 & A;

assign	m3 = B & A;

assign	SYNTHESIZED_WIRE_5 =  ~A;

assign	SYNTHESIZED_WIRE_4 =  ~B;


endmodule
