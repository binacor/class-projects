// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Wed Mar 08 00:27:50 2017"

module in0001(
	n
);


output wire	[15:0] n;

wire	[15:0] n_ALTERA_SYNTHESIZED;






assign	n = n_ALTERA_SYNTHESIZED;
assign	n_ALTERA_SYNTHESIZED[15] = 0;
assign	n_ALTERA_SYNTHESIZED[0] = 1;
assign	n_ALTERA_SYNTHESIZED[14] = 0;
assign	n_ALTERA_SYNTHESIZED[13] = 0;
assign	n_ALTERA_SYNTHESIZED[12] = 0;
assign	n_ALTERA_SYNTHESIZED[11] = 0;
assign	n_ALTERA_SYNTHESIZED[10] = 0;
assign	n_ALTERA_SYNTHESIZED[9] = 0;
assign	n_ALTERA_SYNTHESIZED[8] = 0;
assign	n_ALTERA_SYNTHESIZED[7] = 0;
assign	n_ALTERA_SYNTHESIZED[6] = 0;
assign	n_ALTERA_SYNTHESIZED[5] = 0;
assign	n_ALTERA_SYNTHESIZED[4] = 0;
assign	n_ALTERA_SYNTHESIZED[3] = 0;
assign	n_ALTERA_SYNTHESIZED[2] = 0;
assign	n_ALTERA_SYNTHESIZED[1] = 0;

endmodule
